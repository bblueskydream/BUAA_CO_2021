`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:11:28 11/10/2021 
// Design Name: 
// Module Name:    practice 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module practice(
	input [31:0] in,
	output out
    );
	 reg [31:0] n;
	always@(*)begin
		integer i = 0;
		for (i=0;i<32;i=i+1)begin
		end
	end
	
	always@(*)begin
		n = in;
	end
endmodule
